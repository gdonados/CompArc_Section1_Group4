module or64 (A, B, C);
input [63:0] A, B;  //data inputs
output [63:0] C; //data outputs

C=A|B;

endmodule
