module adderLookAhead64 (A, B, carry, out);
	input [63:0] A, B;
	input carry;
	output [63:0] out;
	
//design a 3-stage carry look-ahead adder 
wire g0, g1, g2, g3, g4


endmodule

//1bit adder
